module chip8

struct Input {
pub mut:
	keys []byte
}

pub fn initialize_input() &Input {
	return &Input{
		keys: []byte{
			len: 16,
			init: 0
		}
	}
}